'timescale 1ns/1ps

module fsm_tb;
    
    reg clk;
    reg reset;
    reg x;
    wire z;


    